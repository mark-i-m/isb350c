`timescale 1ps/1ps

// A toy implementation of the ISB (Jain and Lin, MICRO14).

module isb(input clk); // TODO insert ISB here

endmodule
