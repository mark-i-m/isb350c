`timescale 1ps/1ps

// This is the dispatcher logic. It is mostly a big block
// of combinational logic that was left in its own file.
//
// Inputs:
// CDB
// IB
//
// Outputs:
// ib_flush?
// branch_taken?/branch_target
// REGS
//  - which regs to update
//  - how to update them
// RSs
//  - which RSs to update
//  - what are the values

module dispatch(); //TODO: stuff here

endmodule
